module johnsoncounter( out,reset,clk);
input clk,reset;
output [3:0] out;
reg [3:0] q;
always @(posedge clk)
begin
if(reset)
q=4'd0;
else
begin
q[3]<=q[2];
q[2]<=q[1];
q[1]<=q[0];
q[0]<=(~q[3]);
end

end

assign out=q;

endmodule
