module alu_tb();
reg [3:0]a,b;
reg[3:0]sel;
wire [3:0]y;
wire [7:0]x;
alu dut(a,b,sel,y,x);
initial
begin
sel=4'b0000;a=4'b1010; b=4'b0101;
#5; sel=4'b0001;a=4'b1010; b=4'b0101;
#5; sel=4'b0010;a=4'b1010; b=4'b0101;
#5; sel=4'b0011;a=4'b1010; b=4'b0101;
#5; sel=4'b0100;a=4'b1010; b=4'b0101;
#5; sel=4'b0101;a=4'b1010; b=4'b0101;
#5; sel=4'b0110;a=4'b1010; b=4'b0101;
#5; sel=4'b0111;a=4'b1010; b=4'b0101;
#5; sel=4'b1000;a=4'b1010; b=4'b0101;
#5; sel=4'b1001;a=4'b1010; b=4'b0101;
#5; sel=4'b1010;a=4'b1010; b=4'b0101;
#5; sel=4'b1011;a=4'b1010; b=4'b0101;
#5; sel=4'b1100;a=4'b1010; b=4'b0101;
#5; sel=4'b1101;a=4'b1010; b=4'b0101;
#5; sel=4'b1110;a=4'b1010; b=4'b0101;
#5; sel=4'b1111;a=4'b1010; b=4'b0101;
end

endmodule
