

module decoder3to8(input a,b,cin,
                   output reg[7:0]y
               );


always @(*)
begin
case({a,b,cin})
3'b000:y=8'b00000001;
3'b001:y=8'b00000010;
3'b010:y=8'b00000100;
3'b011:y=8'b00001000;
3'b100:y=8'b00010000;
3'b101:y=8'b00100000;
3'b110:y=8'b01000000;
3'b111:y=8'b10000000;
default:y=8'b00000000;
endcase
end
endmodule


module fuladderwith_decod( 
                           input a,b,cin,
                           
                           output sum,carry
                      
                         );
wire [7:0]w;

decoder3to8 d1(.a(a),.b(b),.cin(cin),.y(w)); 

or o1(sum,w[1],w[2],w[4],w[7]);
or o2(carry,w[3],w[5],w[6],w[7]);
endmodule














